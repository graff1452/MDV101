module register (
    input wire [15:0] d_in,
    input wire reset,
    input wire clk,
    input wire en,
    output reg [15:0] d_out
);

    always @(posedge clk) 
    
endmodule